magic
tech gf180mcuD
magscale 1 5
timestamp 1700650874
<< obsm1 >>
rect 672 855 199304 198382
<< metal2 >>
rect 15904 0 15960 400
rect 16464 0 16520 400
rect 17024 0 17080 400
rect 17584 0 17640 400
rect 18144 0 18200 400
rect 18704 0 18760 400
rect 19264 0 19320 400
rect 19824 0 19880 400
rect 20384 0 20440 400
rect 20944 0 21000 400
rect 21504 0 21560 400
rect 22064 0 22120 400
rect 22624 0 22680 400
rect 23184 0 23240 400
rect 23744 0 23800 400
rect 24304 0 24360 400
rect 24864 0 24920 400
rect 25424 0 25480 400
rect 25984 0 26040 400
rect 26544 0 26600 400
rect 27104 0 27160 400
rect 27664 0 27720 400
rect 28224 0 28280 400
rect 28784 0 28840 400
rect 29344 0 29400 400
rect 29904 0 29960 400
rect 30464 0 30520 400
rect 31024 0 31080 400
rect 31584 0 31640 400
rect 32144 0 32200 400
rect 32704 0 32760 400
rect 33264 0 33320 400
rect 33824 0 33880 400
rect 34384 0 34440 400
rect 34944 0 35000 400
rect 35504 0 35560 400
rect 36064 0 36120 400
rect 36624 0 36680 400
rect 37184 0 37240 400
rect 37744 0 37800 400
rect 38304 0 38360 400
rect 38864 0 38920 400
rect 39424 0 39480 400
rect 39984 0 40040 400
rect 40544 0 40600 400
rect 41104 0 41160 400
rect 41664 0 41720 400
rect 42224 0 42280 400
rect 42784 0 42840 400
rect 43344 0 43400 400
rect 43904 0 43960 400
rect 44464 0 44520 400
rect 45024 0 45080 400
rect 45584 0 45640 400
rect 46144 0 46200 400
rect 46704 0 46760 400
rect 47264 0 47320 400
rect 47824 0 47880 400
rect 48384 0 48440 400
rect 48944 0 49000 400
rect 49504 0 49560 400
rect 50064 0 50120 400
rect 50624 0 50680 400
rect 51184 0 51240 400
rect 51744 0 51800 400
rect 52304 0 52360 400
rect 52864 0 52920 400
rect 53424 0 53480 400
rect 53984 0 54040 400
rect 54544 0 54600 400
rect 55104 0 55160 400
rect 55664 0 55720 400
rect 56224 0 56280 400
rect 56784 0 56840 400
rect 57344 0 57400 400
rect 57904 0 57960 400
rect 58464 0 58520 400
rect 59024 0 59080 400
rect 59584 0 59640 400
rect 60144 0 60200 400
rect 60704 0 60760 400
rect 61264 0 61320 400
rect 61824 0 61880 400
rect 62384 0 62440 400
rect 62944 0 63000 400
rect 63504 0 63560 400
rect 64064 0 64120 400
rect 64624 0 64680 400
rect 65184 0 65240 400
rect 65744 0 65800 400
rect 66304 0 66360 400
rect 66864 0 66920 400
rect 67424 0 67480 400
rect 67984 0 68040 400
rect 68544 0 68600 400
rect 69104 0 69160 400
rect 69664 0 69720 400
rect 70224 0 70280 400
rect 70784 0 70840 400
rect 71344 0 71400 400
rect 71904 0 71960 400
rect 72464 0 72520 400
rect 73024 0 73080 400
rect 73584 0 73640 400
rect 74144 0 74200 400
rect 74704 0 74760 400
rect 75264 0 75320 400
rect 75824 0 75880 400
rect 76384 0 76440 400
rect 76944 0 77000 400
rect 77504 0 77560 400
rect 78064 0 78120 400
rect 78624 0 78680 400
rect 79184 0 79240 400
rect 79744 0 79800 400
rect 80304 0 80360 400
rect 80864 0 80920 400
rect 81424 0 81480 400
rect 81984 0 82040 400
rect 82544 0 82600 400
rect 83104 0 83160 400
rect 83664 0 83720 400
rect 84224 0 84280 400
rect 84784 0 84840 400
rect 85344 0 85400 400
rect 85904 0 85960 400
rect 86464 0 86520 400
rect 87024 0 87080 400
rect 87584 0 87640 400
rect 88144 0 88200 400
rect 88704 0 88760 400
rect 89264 0 89320 400
rect 89824 0 89880 400
rect 90384 0 90440 400
rect 90944 0 91000 400
rect 91504 0 91560 400
rect 92064 0 92120 400
rect 92624 0 92680 400
rect 93184 0 93240 400
rect 93744 0 93800 400
rect 94304 0 94360 400
rect 94864 0 94920 400
rect 95424 0 95480 400
rect 95984 0 96040 400
rect 96544 0 96600 400
rect 97104 0 97160 400
rect 97664 0 97720 400
rect 98224 0 98280 400
rect 98784 0 98840 400
rect 99344 0 99400 400
rect 99904 0 99960 400
rect 100464 0 100520 400
rect 101024 0 101080 400
rect 101584 0 101640 400
rect 102144 0 102200 400
rect 102704 0 102760 400
rect 103264 0 103320 400
rect 103824 0 103880 400
rect 104384 0 104440 400
rect 104944 0 105000 400
rect 105504 0 105560 400
rect 106064 0 106120 400
rect 106624 0 106680 400
rect 107184 0 107240 400
rect 107744 0 107800 400
rect 108304 0 108360 400
rect 108864 0 108920 400
rect 109424 0 109480 400
rect 109984 0 110040 400
rect 110544 0 110600 400
rect 111104 0 111160 400
rect 111664 0 111720 400
rect 112224 0 112280 400
rect 112784 0 112840 400
rect 113344 0 113400 400
rect 113904 0 113960 400
rect 114464 0 114520 400
rect 115024 0 115080 400
rect 115584 0 115640 400
rect 116144 0 116200 400
rect 116704 0 116760 400
rect 117264 0 117320 400
rect 117824 0 117880 400
rect 118384 0 118440 400
rect 118944 0 119000 400
rect 119504 0 119560 400
rect 120064 0 120120 400
rect 120624 0 120680 400
rect 121184 0 121240 400
rect 121744 0 121800 400
rect 122304 0 122360 400
rect 122864 0 122920 400
rect 123424 0 123480 400
rect 123984 0 124040 400
rect 124544 0 124600 400
rect 125104 0 125160 400
rect 125664 0 125720 400
rect 126224 0 126280 400
rect 126784 0 126840 400
rect 127344 0 127400 400
rect 127904 0 127960 400
rect 128464 0 128520 400
rect 129024 0 129080 400
rect 129584 0 129640 400
rect 130144 0 130200 400
rect 130704 0 130760 400
rect 131264 0 131320 400
rect 131824 0 131880 400
rect 132384 0 132440 400
rect 132944 0 133000 400
rect 133504 0 133560 400
rect 134064 0 134120 400
rect 134624 0 134680 400
rect 135184 0 135240 400
rect 135744 0 135800 400
rect 136304 0 136360 400
rect 136864 0 136920 400
rect 137424 0 137480 400
rect 137984 0 138040 400
rect 138544 0 138600 400
rect 139104 0 139160 400
rect 139664 0 139720 400
rect 140224 0 140280 400
rect 140784 0 140840 400
rect 141344 0 141400 400
rect 141904 0 141960 400
rect 142464 0 142520 400
rect 143024 0 143080 400
rect 143584 0 143640 400
rect 144144 0 144200 400
rect 144704 0 144760 400
rect 145264 0 145320 400
rect 145824 0 145880 400
rect 146384 0 146440 400
rect 146944 0 147000 400
rect 147504 0 147560 400
rect 148064 0 148120 400
rect 148624 0 148680 400
rect 149184 0 149240 400
rect 149744 0 149800 400
rect 150304 0 150360 400
rect 150864 0 150920 400
rect 151424 0 151480 400
rect 151984 0 152040 400
rect 152544 0 152600 400
rect 153104 0 153160 400
rect 153664 0 153720 400
rect 154224 0 154280 400
rect 154784 0 154840 400
rect 155344 0 155400 400
rect 155904 0 155960 400
rect 156464 0 156520 400
rect 157024 0 157080 400
rect 157584 0 157640 400
rect 158144 0 158200 400
rect 158704 0 158760 400
rect 159264 0 159320 400
rect 159824 0 159880 400
rect 160384 0 160440 400
rect 160944 0 161000 400
rect 161504 0 161560 400
rect 162064 0 162120 400
rect 162624 0 162680 400
rect 163184 0 163240 400
rect 163744 0 163800 400
rect 164304 0 164360 400
rect 164864 0 164920 400
rect 165424 0 165480 400
rect 165984 0 166040 400
rect 166544 0 166600 400
rect 167104 0 167160 400
rect 167664 0 167720 400
rect 168224 0 168280 400
rect 168784 0 168840 400
rect 169344 0 169400 400
rect 169904 0 169960 400
rect 170464 0 170520 400
rect 171024 0 171080 400
rect 171584 0 171640 400
rect 172144 0 172200 400
rect 172704 0 172760 400
rect 173264 0 173320 400
rect 173824 0 173880 400
rect 174384 0 174440 400
rect 174944 0 175000 400
rect 175504 0 175560 400
rect 176064 0 176120 400
rect 176624 0 176680 400
rect 177184 0 177240 400
rect 177744 0 177800 400
rect 178304 0 178360 400
rect 178864 0 178920 400
rect 179424 0 179480 400
rect 179984 0 180040 400
rect 180544 0 180600 400
rect 181104 0 181160 400
rect 181664 0 181720 400
rect 182224 0 182280 400
rect 182784 0 182840 400
rect 183344 0 183400 400
rect 183904 0 183960 400
<< obsm2 >>
rect 630 430 199122 198371
rect 630 350 15874 430
rect 15990 350 16434 430
rect 16550 350 16994 430
rect 17110 350 17554 430
rect 17670 350 18114 430
rect 18230 350 18674 430
rect 18790 350 19234 430
rect 19350 350 19794 430
rect 19910 350 20354 430
rect 20470 350 20914 430
rect 21030 350 21474 430
rect 21590 350 22034 430
rect 22150 350 22594 430
rect 22710 350 23154 430
rect 23270 350 23714 430
rect 23830 350 24274 430
rect 24390 350 24834 430
rect 24950 350 25394 430
rect 25510 350 25954 430
rect 26070 350 26514 430
rect 26630 350 27074 430
rect 27190 350 27634 430
rect 27750 350 28194 430
rect 28310 350 28754 430
rect 28870 350 29314 430
rect 29430 350 29874 430
rect 29990 350 30434 430
rect 30550 350 30994 430
rect 31110 350 31554 430
rect 31670 350 32114 430
rect 32230 350 32674 430
rect 32790 350 33234 430
rect 33350 350 33794 430
rect 33910 350 34354 430
rect 34470 350 34914 430
rect 35030 350 35474 430
rect 35590 350 36034 430
rect 36150 350 36594 430
rect 36710 350 37154 430
rect 37270 350 37714 430
rect 37830 350 38274 430
rect 38390 350 38834 430
rect 38950 350 39394 430
rect 39510 350 39954 430
rect 40070 350 40514 430
rect 40630 350 41074 430
rect 41190 350 41634 430
rect 41750 350 42194 430
rect 42310 350 42754 430
rect 42870 350 43314 430
rect 43430 350 43874 430
rect 43990 350 44434 430
rect 44550 350 44994 430
rect 45110 350 45554 430
rect 45670 350 46114 430
rect 46230 350 46674 430
rect 46790 350 47234 430
rect 47350 350 47794 430
rect 47910 350 48354 430
rect 48470 350 48914 430
rect 49030 350 49474 430
rect 49590 350 50034 430
rect 50150 350 50594 430
rect 50710 350 51154 430
rect 51270 350 51714 430
rect 51830 350 52274 430
rect 52390 350 52834 430
rect 52950 350 53394 430
rect 53510 350 53954 430
rect 54070 350 54514 430
rect 54630 350 55074 430
rect 55190 350 55634 430
rect 55750 350 56194 430
rect 56310 350 56754 430
rect 56870 350 57314 430
rect 57430 350 57874 430
rect 57990 350 58434 430
rect 58550 350 58994 430
rect 59110 350 59554 430
rect 59670 350 60114 430
rect 60230 350 60674 430
rect 60790 350 61234 430
rect 61350 350 61794 430
rect 61910 350 62354 430
rect 62470 350 62914 430
rect 63030 350 63474 430
rect 63590 350 64034 430
rect 64150 350 64594 430
rect 64710 350 65154 430
rect 65270 350 65714 430
rect 65830 350 66274 430
rect 66390 350 66834 430
rect 66950 350 67394 430
rect 67510 350 67954 430
rect 68070 350 68514 430
rect 68630 350 69074 430
rect 69190 350 69634 430
rect 69750 350 70194 430
rect 70310 350 70754 430
rect 70870 350 71314 430
rect 71430 350 71874 430
rect 71990 350 72434 430
rect 72550 350 72994 430
rect 73110 350 73554 430
rect 73670 350 74114 430
rect 74230 350 74674 430
rect 74790 350 75234 430
rect 75350 350 75794 430
rect 75910 350 76354 430
rect 76470 350 76914 430
rect 77030 350 77474 430
rect 77590 350 78034 430
rect 78150 350 78594 430
rect 78710 350 79154 430
rect 79270 350 79714 430
rect 79830 350 80274 430
rect 80390 350 80834 430
rect 80950 350 81394 430
rect 81510 350 81954 430
rect 82070 350 82514 430
rect 82630 350 83074 430
rect 83190 350 83634 430
rect 83750 350 84194 430
rect 84310 350 84754 430
rect 84870 350 85314 430
rect 85430 350 85874 430
rect 85990 350 86434 430
rect 86550 350 86994 430
rect 87110 350 87554 430
rect 87670 350 88114 430
rect 88230 350 88674 430
rect 88790 350 89234 430
rect 89350 350 89794 430
rect 89910 350 90354 430
rect 90470 350 90914 430
rect 91030 350 91474 430
rect 91590 350 92034 430
rect 92150 350 92594 430
rect 92710 350 93154 430
rect 93270 350 93714 430
rect 93830 350 94274 430
rect 94390 350 94834 430
rect 94950 350 95394 430
rect 95510 350 95954 430
rect 96070 350 96514 430
rect 96630 350 97074 430
rect 97190 350 97634 430
rect 97750 350 98194 430
rect 98310 350 98754 430
rect 98870 350 99314 430
rect 99430 350 99874 430
rect 99990 350 100434 430
rect 100550 350 100994 430
rect 101110 350 101554 430
rect 101670 350 102114 430
rect 102230 350 102674 430
rect 102790 350 103234 430
rect 103350 350 103794 430
rect 103910 350 104354 430
rect 104470 350 104914 430
rect 105030 350 105474 430
rect 105590 350 106034 430
rect 106150 350 106594 430
rect 106710 350 107154 430
rect 107270 350 107714 430
rect 107830 350 108274 430
rect 108390 350 108834 430
rect 108950 350 109394 430
rect 109510 350 109954 430
rect 110070 350 110514 430
rect 110630 350 111074 430
rect 111190 350 111634 430
rect 111750 350 112194 430
rect 112310 350 112754 430
rect 112870 350 113314 430
rect 113430 350 113874 430
rect 113990 350 114434 430
rect 114550 350 114994 430
rect 115110 350 115554 430
rect 115670 350 116114 430
rect 116230 350 116674 430
rect 116790 350 117234 430
rect 117350 350 117794 430
rect 117910 350 118354 430
rect 118470 350 118914 430
rect 119030 350 119474 430
rect 119590 350 120034 430
rect 120150 350 120594 430
rect 120710 350 121154 430
rect 121270 350 121714 430
rect 121830 350 122274 430
rect 122390 350 122834 430
rect 122950 350 123394 430
rect 123510 350 123954 430
rect 124070 350 124514 430
rect 124630 350 125074 430
rect 125190 350 125634 430
rect 125750 350 126194 430
rect 126310 350 126754 430
rect 126870 350 127314 430
rect 127430 350 127874 430
rect 127990 350 128434 430
rect 128550 350 128994 430
rect 129110 350 129554 430
rect 129670 350 130114 430
rect 130230 350 130674 430
rect 130790 350 131234 430
rect 131350 350 131794 430
rect 131910 350 132354 430
rect 132470 350 132914 430
rect 133030 350 133474 430
rect 133590 350 134034 430
rect 134150 350 134594 430
rect 134710 350 135154 430
rect 135270 350 135714 430
rect 135830 350 136274 430
rect 136390 350 136834 430
rect 136950 350 137394 430
rect 137510 350 137954 430
rect 138070 350 138514 430
rect 138630 350 139074 430
rect 139190 350 139634 430
rect 139750 350 140194 430
rect 140310 350 140754 430
rect 140870 350 141314 430
rect 141430 350 141874 430
rect 141990 350 142434 430
rect 142550 350 142994 430
rect 143110 350 143554 430
rect 143670 350 144114 430
rect 144230 350 144674 430
rect 144790 350 145234 430
rect 145350 350 145794 430
rect 145910 350 146354 430
rect 146470 350 146914 430
rect 147030 350 147474 430
rect 147590 350 148034 430
rect 148150 350 148594 430
rect 148710 350 149154 430
rect 149270 350 149714 430
rect 149830 350 150274 430
rect 150390 350 150834 430
rect 150950 350 151394 430
rect 151510 350 151954 430
rect 152070 350 152514 430
rect 152630 350 153074 430
rect 153190 350 153634 430
rect 153750 350 154194 430
rect 154310 350 154754 430
rect 154870 350 155314 430
rect 155430 350 155874 430
rect 155990 350 156434 430
rect 156550 350 156994 430
rect 157110 350 157554 430
rect 157670 350 158114 430
rect 158230 350 158674 430
rect 158790 350 159234 430
rect 159350 350 159794 430
rect 159910 350 160354 430
rect 160470 350 160914 430
rect 161030 350 161474 430
rect 161590 350 162034 430
rect 162150 350 162594 430
rect 162710 350 163154 430
rect 163270 350 163714 430
rect 163830 350 164274 430
rect 164390 350 164834 430
rect 164950 350 165394 430
rect 165510 350 165954 430
rect 166070 350 166514 430
rect 166630 350 167074 430
rect 167190 350 167634 430
rect 167750 350 168194 430
rect 168310 350 168754 430
rect 168870 350 169314 430
rect 169430 350 169874 430
rect 169990 350 170434 430
rect 170550 350 170994 430
rect 171110 350 171554 430
rect 171670 350 172114 430
rect 172230 350 172674 430
rect 172790 350 173234 430
rect 173350 350 173794 430
rect 173910 350 174354 430
rect 174470 350 174914 430
rect 175030 350 175474 430
rect 175590 350 176034 430
rect 176150 350 176594 430
rect 176710 350 177154 430
rect 177270 350 177714 430
rect 177830 350 178274 430
rect 178390 350 178834 430
rect 178950 350 179394 430
rect 179510 350 179954 430
rect 180070 350 180514 430
rect 180630 350 181074 430
rect 181190 350 181634 430
rect 181750 350 182194 430
rect 182310 350 182754 430
rect 182870 350 183314 430
rect 183430 350 183874 430
rect 183990 350 199122 430
<< metal3 >>
rect 0 195216 400 195272
rect 199600 195216 200000 195272
rect 0 186928 400 186984
rect 199600 186928 200000 186984
rect 0 178640 400 178696
rect 199600 178640 200000 178696
rect 0 170352 400 170408
rect 199600 170352 200000 170408
rect 0 162064 400 162120
rect 199600 162064 200000 162120
rect 0 153776 400 153832
rect 199600 153776 200000 153832
rect 0 145488 400 145544
rect 199600 145488 200000 145544
rect 0 137200 400 137256
rect 199600 137200 200000 137256
rect 0 128912 400 128968
rect 199600 128912 200000 128968
rect 0 120624 400 120680
rect 199600 120624 200000 120680
rect 0 112336 400 112392
rect 199600 112336 200000 112392
rect 0 104048 400 104104
rect 199600 104048 200000 104104
rect 0 95760 400 95816
rect 199600 95760 200000 95816
rect 0 87472 400 87528
rect 199600 87472 200000 87528
rect 0 79184 400 79240
rect 199600 79184 200000 79240
rect 0 70896 400 70952
rect 199600 70896 200000 70952
rect 0 62608 400 62664
rect 199600 62608 200000 62664
rect 0 54320 400 54376
rect 199600 54320 200000 54376
rect 0 46032 400 46088
rect 199600 46032 200000 46088
rect 0 37744 400 37800
rect 199600 37744 200000 37800
rect 0 29456 400 29512
rect 199600 29456 200000 29512
rect 0 21168 400 21224
rect 199600 21168 200000 21224
rect 0 12880 400 12936
rect 199600 12880 200000 12936
rect 0 4592 400 4648
rect 199600 4592 200000 4648
<< obsm3 >>
rect 400 195302 199600 198366
rect 430 195186 199570 195302
rect 400 187014 199600 195186
rect 430 186898 199570 187014
rect 400 178726 199600 186898
rect 430 178610 199570 178726
rect 400 170438 199600 178610
rect 430 170322 199570 170438
rect 400 162150 199600 170322
rect 430 162034 199570 162150
rect 400 153862 199600 162034
rect 430 153746 199570 153862
rect 400 145574 199600 153746
rect 430 145458 199570 145574
rect 400 137286 199600 145458
rect 430 137170 199570 137286
rect 400 128998 199600 137170
rect 430 128882 199570 128998
rect 400 120710 199600 128882
rect 430 120594 199570 120710
rect 400 112422 199600 120594
rect 430 112306 199570 112422
rect 400 104134 199600 112306
rect 430 104018 199570 104134
rect 400 95846 199600 104018
rect 430 95730 199570 95846
rect 400 87558 199600 95730
rect 430 87442 199570 87558
rect 400 79270 199600 87442
rect 430 79154 199570 79270
rect 400 70982 199600 79154
rect 430 70866 199570 70982
rect 400 62694 199600 70866
rect 430 62578 199570 62694
rect 400 54406 199600 62578
rect 430 54290 199570 54406
rect 400 46118 199600 54290
rect 430 46002 199570 46118
rect 400 37830 199600 46002
rect 430 37714 199570 37830
rect 400 29542 199600 37714
rect 430 29426 199570 29542
rect 400 21254 199600 29426
rect 430 21138 199570 21254
rect 400 12966 199600 21138
rect 430 12850 199570 12966
rect 400 4678 199600 12850
rect 430 4562 199570 4678
rect 400 406 199600 4562
<< metal4 >>
rect 2224 1538 2384 198382
rect 9904 1538 10064 198382
rect 17584 1538 17744 198382
rect 25264 1538 25424 198382
rect 32944 1538 33104 198382
rect 40624 1538 40784 198382
rect 48304 1538 48464 198382
rect 55984 1538 56144 198382
rect 63664 1538 63824 198382
rect 71344 1538 71504 198382
rect 79024 1538 79184 198382
rect 86704 1538 86864 198382
rect 94384 1538 94544 198382
rect 102064 1538 102224 198382
rect 109744 1538 109904 198382
rect 117424 1538 117584 198382
rect 125104 1538 125264 198382
rect 132784 1538 132944 198382
rect 140464 1538 140624 198382
rect 148144 1538 148304 198382
rect 155824 1538 155984 198382
rect 163504 1538 163664 198382
rect 171184 1538 171344 198382
rect 178864 1538 179024 198382
rect 186544 1538 186704 198382
rect 194224 1538 194384 198382
<< obsm4 >>
rect 2926 1508 9874 179023
rect 10094 1508 17554 179023
rect 17774 1508 25234 179023
rect 25454 1508 32914 179023
rect 33134 1508 40594 179023
rect 40814 1508 48274 179023
rect 48494 1508 55954 179023
rect 56174 1508 63634 179023
rect 63854 1508 71314 179023
rect 71534 1508 78994 179023
rect 79214 1508 86674 179023
rect 86894 1508 94354 179023
rect 94574 1508 102034 179023
rect 102254 1508 109714 179023
rect 109934 1508 117394 179023
rect 117614 1508 125074 179023
rect 125294 1508 126434 179023
rect 2926 569 126434 1508
<< labels >>
rlabel metal3 s 199600 4592 200000 4648 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 145488 400 145544 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 120624 400 120680 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 95760 400 95816 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 70896 400 70952 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 46032 400 46088 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 21168 400 21224 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 199600 29456 200000 29512 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 199600 54320 200000 54376 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 199600 79184 200000 79240 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 199600 104048 200000 104104 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 199600 128912 200000 128968 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 199600 153776 200000 153832 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 199600 178640 200000 178696 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 195216 400 195272 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 170352 400 170408 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 199600 21168 200000 21224 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 128912 400 128968 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 104048 400 104104 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 79184 400 79240 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 54320 400 54376 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 29456 400 29512 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4592 400 4648 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 199600 46032 200000 46088 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 199600 70896 200000 70952 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 199600 95760 200000 95816 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 199600 120624 200000 120680 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 199600 145488 200000 145544 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 199600 170352 200000 170408 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 199600 195216 200000 195272 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 178640 400 178696 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 153776 400 153832 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 199600 12880 200000 12936 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 137200 400 137256 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 112336 400 112392 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 87472 400 87528 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 62608 400 62664 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 37744 400 37800 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 12880 400 12936 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 199600 37744 200000 37800 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 199600 62608 200000 62664 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 199600 87472 200000 87528 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 199600 112336 200000 112392 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 199600 137200 200000 137256 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 199600 162064 200000 162120 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 199600 186928 200000 186984 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 186928 400 186984 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 162064 400 162120 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 182784 0 182840 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 183344 0 183400 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 183904 0 183960 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 75264 0 75320 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 92064 0 92120 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 93744 0 93800 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 95424 0 95480 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 97104 0 97160 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 98784 0 98840 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 100464 0 100520 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 102144 0 102200 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 103824 0 103880 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 105504 0 105560 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 107184 0 107240 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 76944 0 77000 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 108864 0 108920 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 110544 0 110600 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 112224 0 112280 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 113904 0 113960 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 115584 0 115640 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 117264 0 117320 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 118944 0 119000 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 120624 0 120680 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 122304 0 122360 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 123984 0 124040 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 78624 0 78680 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 125664 0 125720 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 127344 0 127400 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 129024 0 129080 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 130704 0 130760 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 132384 0 132440 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 134064 0 134120 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 135744 0 135800 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 137424 0 137480 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 139104 0 139160 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 140784 0 140840 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 80304 0 80360 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 142464 0 142520 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 144144 0 144200 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 145824 0 145880 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 147504 0 147560 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 149184 0 149240 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 150864 0 150920 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 152544 0 152600 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 154224 0 154280 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 155904 0 155960 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 157584 0 157640 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 81984 0 82040 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 159264 0 159320 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 160944 0 161000 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 162624 0 162680 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 164304 0 164360 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 165984 0 166040 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 167664 0 167720 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 169344 0 169400 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 171024 0 171080 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 172704 0 172760 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 174384 0 174440 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 83664 0 83720 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 176064 0 176120 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 177744 0 177800 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 179424 0 179480 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 181104 0 181160 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 85344 0 85400 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 88704 0 88760 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 90384 0 90440 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 75824 0 75880 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 92624 0 92680 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 94304 0 94360 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 95984 0 96040 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 97664 0 97720 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 99344 0 99400 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 101024 0 101080 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 102704 0 102760 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 104384 0 104440 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 106064 0 106120 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 107744 0 107800 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 77504 0 77560 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 111104 0 111160 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 112784 0 112840 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 114464 0 114520 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 116144 0 116200 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 117824 0 117880 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 119504 0 119560 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 121184 0 121240 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 122864 0 122920 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 124544 0 124600 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 79184 0 79240 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 126224 0 126280 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 127904 0 127960 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 129584 0 129640 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 131264 0 131320 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 132944 0 133000 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 134624 0 134680 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 136304 0 136360 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 137984 0 138040 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 139664 0 139720 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 141344 0 141400 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 80864 0 80920 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 143024 0 143080 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 144704 0 144760 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 146384 0 146440 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 148064 0 148120 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 149744 0 149800 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 151424 0 151480 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 153104 0 153160 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 154784 0 154840 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 156464 0 156520 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 158144 0 158200 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 82544 0 82600 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 159824 0 159880 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 161504 0 161560 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 163184 0 163240 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 164864 0 164920 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 166544 0 166600 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 168224 0 168280 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 169904 0 169960 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 171584 0 171640 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 173264 0 173320 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 174944 0 175000 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 84224 0 84280 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 176624 0 176680 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 178304 0 178360 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 179984 0 180040 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 181664 0 181720 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 85904 0 85960 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 87584 0 87640 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 89264 0 89320 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 90944 0 91000 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 76384 0 76440 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 93184 0 93240 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 94864 0 94920 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 96544 0 96600 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 98224 0 98280 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 99904 0 99960 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 101584 0 101640 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 103264 0 103320 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 104944 0 105000 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 106624 0 106680 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 108304 0 108360 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 78064 0 78120 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 109984 0 110040 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 111664 0 111720 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 113344 0 113400 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 115024 0 115080 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 116704 0 116760 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 118384 0 118440 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 120064 0 120120 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 121744 0 121800 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 123424 0 123480 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 125104 0 125160 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 79744 0 79800 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 126784 0 126840 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 128464 0 128520 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 130144 0 130200 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 131824 0 131880 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 133504 0 133560 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 135184 0 135240 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 136864 0 136920 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 138544 0 138600 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 140224 0 140280 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 141904 0 141960 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 81424 0 81480 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 143584 0 143640 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 145264 0 145320 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 146944 0 147000 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 148624 0 148680 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 150304 0 150360 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 151984 0 152040 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 153664 0 153720 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 155344 0 155400 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 157024 0 157080 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 158704 0 158760 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 83104 0 83160 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 160384 0 160440 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 162064 0 162120 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 163744 0 163800 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 165424 0 165480 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 167104 0 167160 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 168784 0 168840 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 170464 0 170520 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 172144 0 172200 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 173824 0 173880 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 175504 0 175560 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 84784 0 84840 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 177184 0 177240 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 178864 0 178920 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 180544 0 180600 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 182224 0 182280 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 86464 0 86520 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 88144 0 88200 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 89824 0 89880 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 91504 0 91560 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 198382 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 198382 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 15904 0 15960 400 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 16464 0 16520 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 17024 0 17080 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 19264 0 19320 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 39984 0 40040 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 41664 0 41720 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 43344 0 43400 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 45024 0 45080 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 48384 0 48440 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 50064 0 50120 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 53424 0 53480 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 55104 0 55160 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 56784 0 56840 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 58464 0 58520 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 61824 0 61880 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 63504 0 63560 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 65184 0 65240 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 68544 0 68600 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 70224 0 70280 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 23744 0 23800 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 71904 0 71960 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 29904 0 29960 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 36624 0 36680 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 38864 0 38920 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 45584 0 45640 400 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 50624 0 50680 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 52304 0 52360 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 57344 0 57400 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 62384 0 62440 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 64064 0 64120 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 65744 0 65800 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 69104 0 69160 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 72464 0 72520 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 74144 0 74200 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 30464 0 30520 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 33824 0 33880 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 37184 0 37240 400 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 39424 0 39480 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 41104 0 41160 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 42784 0 42840 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 44464 0 44520 400 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 46144 0 46200 400 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 47824 0 47880 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 49504 0 49560 400 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 51184 0 51240 400 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 52864 0 52920 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 54544 0 54600 400 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 56224 0 56280 400 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 57904 0 57960 400 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 59584 0 59640 400 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 61264 0 61320 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 62944 0 63000 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 64624 0 64680 400 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 66304 0 66360 400 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 67984 0 68040 400 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 69664 0 69720 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 71344 0 71400 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 24864 0 24920 400 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 73024 0 73080 400 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 74704 0 74760 400 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 27104 0 27160 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 29344 0 29400 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 31024 0 31080 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 32704 0 32760 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 34384 0 34440 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 36064 0 36120 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 37744 0 37800 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 20944 0 21000 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 23184 0 23240 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 25424 0 25480 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 27664 0 27720 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 60063814
string GDS_FILE /home/shahid/Desktop/test123/caravel_user_project/openlane/user_proj_example/runs/23_11_22_14_18/results/signoff/user_proj_example.magic.gds
string GDS_START 609120
<< end >>

